class ex4_agent extends uvm_component;
  //UVM Factory Registration Macro
  `uvm_component_utils(ex4_agent)