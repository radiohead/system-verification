`include "uvm_macros.svh"

package ex1_pkg;
  import uvm_pkg::*;

  `include "ex1_driver.svh"
  `include "ex1_env.svh"
endpackage: ex1_pkg